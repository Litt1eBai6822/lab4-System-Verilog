module vga_controller (
    input logic clk,
    input logic rst,
    output logic hsync,
    output logic vsync,
    output logic [3:0] r,
    output logic [3:0] g,
    output logic [3:0] b
);

// Implementation of VGA controller here

endmodule